// 2023-12/30
// Verilog表达式

// 表达式
a^b; // a异或b
address[9:0] + 10'b01; //地址累加
flag1 && flag2; //逻辑与


// 操作数
// 操作数可以是任意的数据类型，只是某些特定的语法结构要求使用特定类型的操作数。
// 操作数可以为常数，整数，实数，线网，寄存器，时间，位选，域选，存储器及函数调用等。
// always块里赋值对象不能是wire型
// Example:
module test;


//实数
real a, b, c;
c = a + b ;


//寄存器
reg  [3:0]       cprmu_1, cprmu_2 ;
always @(posedge clk) begin  // 时钟沿上升即运算
        cprmu_2 = cprmu_1 ^ cprmu_2 ;
end
         
//函数
reg  flag1 ;
flag = calculate_result(A, B);
 
//非法操作数
reg [3:0]         res;
wire [3:0]        temp;
always@ （*）begin
    res    = cprmu_2 – cprmu_1 ;
    //temp = cprmu_2 – cprmu_1 ; //不合法，always块里赋值对象不能是wire型
end

endmodule


// 双目运算符中，如果有一个操作数是x, 则结果也会是x


// 负数的表示
// 在表示位宽的数字前加符号 例如：
-4 = -4b'0100


// 按位操作符
// 包括：取反（~），与（&），或（|），异或（^），同或（~^）。
// 例如：
A = 4'b0101 ;
B = 4'b1001 ;
C = 4'bx010 ;
    
~A        //4'b1010
A & B     //4'b0001
A | B     //4'b1101
A^B       //4'b1100
A ~^ B    //4'b0011
B | C     //4'b1011
B&C       //4'bx000


// 规约操作符 &, ~&, |, ~| 只有一个操作数， 是按照位数进行运算, 结果是1位
A = 4'b1010 ;
&A ;      //结果为 1 & 0 & 1 & 0 = 1'b0，可用来判断变量A是否全1
~|A ;     //结果为 ~(1 | 0 | 1 | 0) = 1'b0, 可用来判断变量A是否为全0
^A ;      //结果为 1 ^ 0 ^ 1 ^ 0 = 1'b0


// 拼接操作符 {, }
// 拼接符操作数必须指定位宽，常数的话也需要指定位宽。例如：

A = 4'b1010 ;
B = 1'b1 ;
Y1 = {B, A[3:2], A[0], 4'h3 };  //结果为Y1='b1100_0011
Y2 = {4{B}, 3'd4};  //结果为 Y2=7'b111_1100
Y3 = {32{1'b0}};  //结果为 Y3=32h0，常用作寄存器初始化时匹配位宽的赋初值




















